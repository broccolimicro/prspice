* This setting performs a sophisticated path search to all
* feasible power supplies associated with every element and
* node. It detects PWL/PULSE power supplies and internal power
* supply nodes and sets correct voltage supply values.
.param HSIMVDD=1.0v
.param HSIMALLOWEDDV=0.001v
.param HSIMVHTH=0.7v
.param HSIMVLTH=0.3v

* Valid values are: fsdb (the default), wdf, vpd, nassda, out, and alint.
.param HSIMOUTPUT="fsdb&alint"
.param HSIMOUTPUTFLUSH=1n

* Report the average capacitance of the whole circuit
.param HSIMNODECAP="*"

* Lists model statistics in the log file.
.param HSIMMODELSTAT=1

* This setting precisely models and simulates the coupling effects
* between each pair of gate/drain/source/bulk terminals for each
* MOSFET
.param HSIMSPICE=2
.param HSIMB4REMOVE=0
.param HSIMSTEADYCURRENT=1n

* different time stepsizes are selected in
* different subcircuits, such that a smaller time step is
* selected for subcircuits with faster transient activities,
* while a larger time step is selected for subcircuits with
* slow transient activities. This speed-up in multirate step
* selection is achieved by reducing the total number of time
* steps.
.param HSIMSPEED=1
.param HSIMANALOG=2

* Performs a sanity check to identify potential forward bias conditions in
* MOSFET parasitic diodes.
.param HSIMCHECKMOSBULK=1

* Calculates the dc current of MOSFET diodes.
.param HSIMDIODECURRENT=1

* Uses the HSIM proprietary iteration scheme, which
* balances accuracy and performance.
.param HSIMITERMODE=1

* Calculates the static gate leakage currents and the substrate current.
* Includes both the static gate leakage currents and the
* substrate current in the calculation.
.param HSIMIGISUB=1

.param HSIMRISE=30ps
.param HSIMFALL=30ps
